--
-- Inferrable Synchronous SRAM for Leonardo synthesis, no write through!
--
-- Version : 0236
--
-- Copyright (c) 2002 Daniel Wallner (jesus@opencores.org)
--
-- All rights reserved
--
-- Redistribution and use in source and synthezised forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- Redistributions of source code must retain the above copyright notice,
-- this list of conditions and the following disclaimer.
--
-- Redistributions in synthesized form must reproduce the above copyright
-- notice, this list of conditions and the following disclaimer in the
-- documentation and/or other materials provided with the distribution.
--
-- Neither the name of the author nor the names of other contributors may
-- be used to endorse or promote products derived from this software without
-- specific prior written permission.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
--
-- Please report bugs to the author, but before you do so, please
-- make sure that this is not a derivative work and that
-- you have the latest version of this file.
--
-- The latest version of this file can be found at:
--    http://www.opencores.org/cvsweb.shtml/t51/
--
-- Limitations :
--
-- File history :
--

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity $$$ENTITY$$$ is
    generic(
        AddrWidth    : integer := 16;
        DataWidth    : integer := 8
    );
    port(
        Clk         : in std_logic;
        CE_n        : in std_logic;
        WE_n        : in std_logic;
        A           : in std_logic_vector(AddrWidth - 1 downto 0);
        DIn         : in std_logic_vector(DataWidth - 1 downto 0);
        DOut        : out std_logic_vector(DataWidth - 1 downto 0)
    );
end $$$ENTITY$$$;

architecture behaviour of $$$ENTITY$$$ is

    type Memory_Image is array (natural range <>) of std_logic_vector(DataWidth - 1 downto 0);
    signal MemArray: Memory_Image(0 to 2 ** AddrWidth - 1) := (
$$$CONTENT$$$,
        others => X"00"
    );
--    signal    A_r: std_logic_vector(AddrWidth - 1 downto 0);

begin

    process (CE_n, WE_n)
    begin
        if CE_n'event or WE_n'event then
            if CE_n = '0' and WE_n = '1' then
                assert not is_x(A) report "Read from X address" severity FAILURE;
                DOut <= MemArray(to_integer(unsigned(A(AddrWidth - 1 downto 0))));
            end if;
            if CE_n = '0' and WE_n'event and WE_n = '1' then -- we right on the rising edge of CLK, not on the falling one
                assert not is_x(A) report "Write to X address" severity FAILURE;
                assert not is_x(DIn) report "Write X data" severity FAILURE;
                MemArray(to_integer(unsigned(A))) <= DIn;
            end if;
--            A_r <= A;
        end if;
    end process;

end;
